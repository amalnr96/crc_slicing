`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 14.05.2023 23:30:17
// Design Name: 
// Module Name: slicing_by8
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module slicing_by8(

input wire[63:0] data_i, 
input wire[31:0] old_crc_i, 
input wire clk_i, 
input wire rst_i, 
output reg [31:0] new_crc_o

    );
 logic [31:0] crctable0[256]= {32'h00000000,32'h77073096,32'hee0e612c,32'h990951ba,32'h076dc419,32'h706af48f,32'he963a535,32'h9e6495a3,
                               32'h0edb8832,32'h79dcb8a4,32'he0d5e91e,32'h97d2d988,32'h09b64c2b,32'h7eb17cbd,32'he7b82d07,32'h90bf1d91,
                               32'h1db71064,32'h6ab020f2,32'hf3b97148,32'h84be41de,32'h1adad47d,32'h6ddde4eb,32'hf4d4b551,32'h83d385c7,
                               32'h136c9856,32'h646ba8c0,32'hfd62f97a,32'h8a65c9ec,32'h14015c4f,32'h63066cd9,32'hfa0f3d63,32'h8d080df5,
                               32'h3b6e20c8,32'h4c69105e,32'hd56041e4,32'ha2677172,32'h3c03e4d1,32'h4b04d447,32'hd20d85fd,32'ha50ab56b,
                               32'h35b5a8fa,32'h42b2986c,32'hdbbbc9d6,32'hacbcf940,32'h32d86ce3,32'h45df5c75,32'hdcd60dcf,32'habd13d59,
                               32'h26d930ac,32'h51de003a,32'hc8d75180,32'hbfd06116,32'h21b4f4b5,32'h56b3c423,32'hcfba9599,32'hb8bda50f,
                               32'h2802b89e,32'h5f058808,32'hc60cd9b2,32'hb10be924,32'h2f6f7c87,32'h58684c11,32'hc1611dab,32'hb6662d3d,
                               32'h76dc4190,32'h01db7106,32'h98d220bc,32'hefd5102a,32'h71b18589,32'h06b6b51f,32'h9fbfe4a5,32'he8b8d433,
                               32'h7807c9a2,32'h0f00f934,32'h9609a88e,32'he10e9818,32'h7f6a0dbb,32'h086d3d2d,32'h91646c97,32'he6635c01,
                               32'h6b6b51f4,32'h1c6c6162,32'h856530d8,32'hf262004e,32'h6c0695ed,32'h1b01a57b,32'h8208f4c1,32'hf50fc457,
                               32'h65b0d9c6,32'h12b7e950,32'h8bbeb8ea,32'hfcb9887c,32'h62dd1ddf,32'h15da2d49,32'h8cd37cf3,32'hfbd44c65,
                               32'h4db26158,32'h3ab551ce,32'ha3bc0074,32'hd4bb30e2,32'h4adfa541,32'h3dd895d7,32'ha4d1c46d,32'hd3d6f4fb,
                               32'h4369e96a,32'h346ed9fc,32'had678846,32'hda60b8d0,32'h44042d73,32'h33031de5,32'haa0a4c5f,32'hdd0d7cc9,
                               32'h5005713c,32'h270241aa,32'hbe0b1010,32'hc90c2086,32'h5768b525,32'h206f85b3,32'hb966d409,32'hce61e49f,
                               32'h5edef90e,32'h29d9c998,32'hb0d09822,32'hc7d7a8b4,32'h59b33d17,32'h2eb40d81,32'hb7bd5c3b,32'hc0ba6cad,
                               32'hedb88320,32'h9abfb3b6,32'h03b6e20c,32'h74b1d29a,32'head54739,32'h9dd277af,32'h04db2615,32'h73dc1683,
                               32'he3630b12,32'h94643b84,32'h0d6d6a3e,32'h7a6a5aa8,32'he40ecf0b,32'h9309ff9d,32'h0a00ae27,32'h7d079eb1,
                               32'hf00f9344,32'h8708a3d2,32'h1e01f268,32'h6906c2fe,32'hf762575d,32'h806567cb,32'h196c3671,32'h6e6b06e7,
                               32'hfed41b76,32'h89d32be0,32'h10da7a5a,32'h67dd4acc,32'hf9b9df6f,32'h8ebeeff9,32'h17b7be43,32'h60b08ed5,
                               32'hd6d6a3e8,32'ha1d1937e,32'h38d8c2c4,32'h4fdff252,32'hd1bb67f1,32'ha6bc5767,32'h3fb506dd,32'h48b2364b,
                               32'hd80d2bda,32'haf0a1b4c,32'h36034af6,32'h41047a60,32'hdf60efc3,32'ha867df55,32'h316e8eef,32'h4669be79,
                               32'hcb61b38c,32'hbc66831a,32'h256fd2a0,32'h5268e236,32'hcc0c7795,32'hbb0b4703,32'h220216b9,32'h5505262f,
                               32'hc5ba3bbe,32'hb2bd0b28,32'h2bb45a92,32'h5cb36a04,32'hc2d7ffa7,32'hb5d0cf31,32'h2cd99e8b,32'h5bdeae1d,
                               32'h9b64c2b0,32'hec63f226,32'h756aa39c,32'h026d930a,32'h9c0906a9,32'heb0e363f,32'h72076785,32'h05005713,
                               32'h95bf4a82,32'he2b87a14,32'h7bb12bae,32'h0cb61b38,32'h92d28e9b,32'he5d5be0d,32'h7cdcefb7,32'h0bdbdf21,
                               32'h86d3d2d4,32'hf1d4e242,32'h68ddb3f8,32'h1fda836e,32'h81be16cd,32'hf6b9265b,32'h6fb077e1,32'h18b74777,
                               32'h88085ae6,32'hff0f6a70,32'h66063bca,32'h11010b5c,32'h8f659eff,32'hf862ae69,32'h616bffd3,32'h166ccf45,
                               32'ha00ae278,32'hd70dd2ee,32'h4e048354,32'h3903b3c2,32'ha7672661,32'hd06016f7,32'h4969474d,32'h3e6e77db,
                               32'haed16a4a,32'hd9d65adc,32'h40df0b66,32'h37d83bf0,32'ha9bcae53,32'hdebb9ec5,32'h47b2cf7f,32'h30b5ffe9,
                               32'hbdbdf21c,32'hcabac28a,32'h53b39330,32'h24b4a3a6,32'hbad03605,32'hcdd70693,32'h54de5729,32'h23d967bf,
                               32'hb3667a2e,32'hc4614ab8,32'h5d681b02,32'h2a6f2b94,32'hb40bbe37,32'hc30c8ea1,32'h5a05df1b,32'h001c09bc};

 logic [31:0] crctable1[256]= { 32'h00000000,32'h191B3141,32'h32366282,32'h2B2D53C3,32'h646CC504,32'h7D77F445,32'h565AA786,32'h4F4196C7,
    32'hC8D98A08,32'hD1C2BB49,32'hFAEFE88A,32'hE3F4D9CB,32'hACB54F0C,32'hB5AE7E4D,32'h9E832D8E,32'h87981CCF,
    32'h4AC21251,32'h53D92310,32'h78F470D3,32'h61EF4192,32'h2EAED755,32'h37B5E614,32'h1C98B5D7,32'h05838496,
    32'h821B9859,32'h9B00A918,32'hB02DFADB,32'hA936CB9A,32'hE6775D5D,32'hFF6C6C1C,32'hD4413FDF,32'hCD5A0E9E,
    32'h958424A2,32'h8C9F15E3,32'hA7B24620,32'hBEA97761,32'hF1E8E1A6,32'hE8F3D0E7,32'hC3DE8324,32'hDAC5B265,
    32'h5D5DAEAA,32'h44469FEB,32'h6F6BCC28,32'h7670FD69,32'h39316BAE,32'h202A5AEF,32'h0B07092C,32'h121C386D,
    32'hDF4636F3,32'hC65D07B2,32'hED705471,32'hF46B6530,32'hBB2AF3F7,32'hA231C2B6,32'h891C9175,32'h9007A034,
    32'h179FBCFB,32'h0E848DBA,32'h25A9DE79,32'h3CB2EF38,32'h73F379FF,32'h6AE848BE,32'h41C51B7D,32'h58DE2A3C,
    32'hF0794F05,32'hE9627E44,32'hC24F2D87,32'hDB541CC6,32'h94158A01,32'h8D0EBB40,32'hA623E883,32'hBF38D9C2,
    32'h38A0C50D,32'h21BBF44C,32'h0A96A78F,32'h138D96CE,32'h5CCC0009,32'h45D73148,32'h6EFA628B,32'h77E153CA,
    32'hBABB5D54,32'hA3A06C15,32'h888D3FD6,32'h91960E97,32'hDED79850,32'hC7CCA911,32'hECE1FAD2,32'hF5FACB93,
    32'h7262D75C,32'h6B79E61D,32'h4054B5DE,32'h594F849F,32'h160E1258,32'h0F152319,32'h243870DA,32'h3D23419B,
    32'h65FD6BA7,32'h7CE65AE6,32'h57CB0925,32'h4ED03864,32'h0191AEA3,32'h188A9FE2,32'h33A7CC21,32'h2ABCFD60,
    32'hAD24E1AF,32'hB43FD0EE,32'h9F12832D,32'h8609B26C,32'hC94824AB,32'hD05315EA,32'hFB7E4629,32'hE2657768,
    32'h2F3F79F6,32'h362448B7,32'h1D091B74,32'h04122A35,32'h4B53BCF2,32'h52488DB3,32'h7965DE70,32'h607EEF31,
    32'hE7E6F3FE,32'hFEFDC2BF,32'hD5D0917C,32'hCCCBA03D,32'h838A36FA,32'h9A9107BB,32'hB1BC5478,32'hA8A76539,
    32'h3B83984B,32'h2298A90A,32'h09B5FAC9,32'h10AECB88,32'h5FEF5D4F,32'h46F46C0E,32'h6DD93FCD,32'h74C20E8C,
    32'hF35A1243,32'hEA412302,32'hC16C70C1,32'hD8774180,32'h9736D747,32'h8E2DE606,32'hA500B5C5,32'hBC1B8484,
    32'h71418A1A,32'h685ABB5B,32'h4377E898,32'h5A6CD9D9,32'h152D4F1E,32'h0C367E5F,32'h271B2D9C,32'h3E001CDD,
    32'hB9980012,32'hA0833153,32'h8BAE6290,32'h92B553D1,32'hDDF4C516,32'hC4EFF457,32'hEFC2A794,32'hF6D996D5,
    32'hAE07BCE9,32'hB71C8DA8,32'h9C31DE6B,32'h852AEF2A,32'hCA6B79ED,32'hD37048AC,32'hF85D1B6F,32'hE1462A2E,
    32'h66DE36E1,32'h7FC507A0,32'h54E85463,32'h4DF36522,32'h02B2F3E5,32'h1BA9C2A4,32'h30849167,32'h299FA026,
    32'hE4C5AEB8,32'hFDDE9FF9,32'hD6F3CC3A,32'hCFE8FD7B,32'h80A96BBC,32'h99B25AFD,32'hB29F093E,32'hAB84387F,
    32'h2C1C24B0,32'h350715F1,32'h1E2A4632,32'h07317773,32'h4870E1B4,32'h516BD0F5,32'h7A468336,32'h635DB277,
    32'hCBFAD74E,32'hD2E1E60F,32'hF9CCB5CC,32'hE0D7848D,32'hAF96124A,32'hB68D230B,32'h9DA070C8,32'h84BB4189,
    32'h03235D46,32'h1A386C07,32'h31153FC4,32'h280E0E85,32'h674F9842,32'h7E54A903,32'h5579FAC0,32'h4C62CB81,
    32'h8138C51F,32'h9823F45E,32'hB30EA79D,32'hAA1596DC,32'hE554001B,32'hFC4F315A,32'hD7626299,32'hCE7953D8,
    32'h49E14F17,32'h50FA7E56,32'h7BD72D95,32'h62CC1CD4,32'h2D8D8A13,32'h3496BB52,32'h1FBBE891,32'h06A0D9D0,
    32'h5E7EF3EC,32'h4765C2AD,32'h6C48916E,32'h7553A02F,32'h3A1236E8,32'h230907A9,32'h0824546A,32'h113F652B,
    32'h96A779E4,32'h8FBC48A5,32'hA4911B66,32'hBD8A2A27,32'hF2CBBCE0,32'hEBD08DA1,32'hC0FDDE62,32'hD9E6EF23,
    32'h14BCE1BD,32'h0DA7D0FC,32'h268A833F,32'h3F91B27E,32'h70D024B9,32'h69CB15F8,32'h42E6463B,32'h5BFD777A,
    32'hDC656BB5,32'hC57E5AF4,32'hEE530937,32'hF7483876,32'hB809AEB1,32'hA1129FF0,32'h8A3FCC33,32'h9324FD72};

 logic [31:0] crctable2[256]= {32'h00000000,32'h01C26A37,32'h0384D46E,32'h0246BE59,32'h0709A8DC,32'h06CBC2EB,32'h048D7CB2,32'h054F1685,
    32'h0E1351B8,32'h0FD13B8F,32'h0D9785D6,32'h0C55EFE1,32'h091AF964,32'h08D89353,32'h0A9E2D0A,32'h0B5C473D,
    32'h1C26A370,32'h1DE4C947,32'h1FA2771E,32'h1E601D29,32'h1B2F0BAC,32'h1AED619B,32'h18ABDFC2,32'h1969B5F5,
    32'h1235F2C8,32'h13F798FF,32'h11B126A6,32'h10734C91,32'h153C5A14,32'h14FE3023,32'h16B88E7A,32'h177AE44D,
    32'h384D46E0,32'h398F2CD7,32'h3BC9928E,32'h3A0BF8B9,32'h3F44EE3C,32'h3E86840B,32'h3CC03A52,32'h3D025065,
    32'h365E1758,32'h379C7D6F,32'h35DAC336,32'h3418A901,32'h3157BF84,32'h3095D5B3,32'h32D36BEA,32'h331101DD,
    32'h246BE590,32'h25A98FA7,32'h27EF31FE,32'h262D5BC9,32'h23624D4C,32'h22A0277B,32'h20E69922,32'h2124F315,
    32'h2A78B428,32'h2BBADE1F,32'h29FC6046,32'h283E0A71,32'h2D711CF4,32'h2CB376C3,32'h2EF5C89A,32'h2F37A2AD,
    32'h709A8DC0,32'h7158E7F7,32'h731E59AE,32'h72DC3399,32'h7793251C,32'h76514F2B,32'h7417F172,32'h75D59B45,
    32'h7E89DC78,32'h7F4BB64F,32'h7D0D0816,32'h7CCF6221,32'h798074A4,32'h78421E93,32'h7A04A0CA,32'h7BC6CAFD,
    32'h6CBC2EB0,32'h6D7E4487,32'h6F38FADE,32'h6EFA90E9,32'h6BB5866C,32'h6A77EC5B,32'h68315202,32'h69F33835,
    32'h62AF7F08,32'h636D153F,32'h612BAB66,32'h60E9C151,32'h65A6D7D4,32'h6464BDE3,32'h662203BA,32'h67E0698D,
    32'h48D7CB20,32'h4915A117,32'h4B531F4E,32'h4A917579,32'h4FDE63FC,32'h4E1C09CB,32'h4C5AB792,32'h4D98DDA5,
    32'h46C49A98,32'h4706F0AF,32'h45404EF6,32'h448224C1,32'h41CD3244,32'h400F5873,32'h4249E62A,32'h438B8C1D,
    32'h54F16850,32'h55330267,32'h5775BC3E,32'h56B7D609,32'h53F8C08C,32'h523AAABB,32'h507C14E2,32'h51BE7ED5,
    32'h5AE239E8,32'h5B2053DF,32'h5966ED86,32'h58A487B1,32'h5DEB9134,32'h5C29FB03,32'h5E6F455A,32'h5FAD2F6D,
    32'hE1351B80,32'hE0F771B7,32'hE2B1CFEE,32'hE373A5D9,32'hE63CB35C,32'hE7FED96B,32'hE5B86732,32'hE47A0D05,
    32'hEF264A38,32'hEEE4200F,32'hECA29E56,32'hED60F461,32'hE82FE2E4,32'hE9ED88D3,32'hEBAB368A,32'hEA695CBD,
    32'hFD13B8F0,32'hFCD1D2C7,32'hFE976C9E,32'hFF5506A9,32'hFA1A102C,32'hFBD87A1B,32'hF99EC442,32'hF85CAE75,
    32'hF300E948,32'hF2C2837F,32'hF0843D26,32'hF1465711,32'hF4094194,32'hF5CB2BA3,32'hF78D95FA,32'hF64FFFCD,
    32'hD9785D60,32'hD8BA3757,32'hDAFC890E,32'hDB3EE339,32'hDE71F5BC,32'hDFB39F8B,32'hDDF521D2,32'hDC374BE5,
    32'hD76B0CD8,32'hD6A966EF,32'hD4EFD8B6,32'hD52DB281,32'hD062A404,32'hD1A0CE33,32'hD3E6706A,32'hD2241A5D,
    32'hC55EFE10,32'hC49C9427,32'hC6DA2A7E,32'hC7184049,32'hC25756CC,32'hC3953CFB,32'hC1D382A2,32'hC011E895,
    32'hCB4DAFA8,32'hCA8FC59F,32'hC8C97BC6,32'hC90B11F1,32'hCC440774,32'hCD866D43,32'hCFC0D31A,32'hCE02B92D,
    32'h91AF9640,32'h906DFC77,32'h922B422E,32'h93E92819,32'h96A63E9C,32'h976454AB,32'h9522EAF2,32'h94E080C5,
    32'h9FBCC7F8,32'h9E7EADCF,32'h9C381396,32'h9DFA79A1,32'h98B56F24,32'h99770513,32'h9B31BB4A,32'h9AF3D17D,
    32'h8D893530,32'h8C4B5F07,32'h8E0DE15E,32'h8FCF8B69,32'h8A809DEC,32'h8B42F7DB,32'h89044982,32'h88C623B5,
    32'h839A6488,32'h82580EBF,32'h801EB0E6,32'h81DCDAD1,32'h8493CC54,32'h8551A663,32'h8717183A,32'h86D5720D,
    32'hA9E2D0A0,32'hA820BA97,32'hAA6604CE,32'hABA46EF9,32'hAEEB787C,32'hAF29124B,32'hAD6FAC12,32'hACADC625,
    32'hA7F18118,32'hA633EB2F,32'hA4755576,32'hA5B73F41,32'hA0F829C4,32'hA13A43F3,32'hA37CFDAA,32'hA2BE979D,
    32'hB5C473D0,32'hB40619E7,32'hB640A7BE,32'hB782CD89,32'hB2CDDB0C,32'hB30FB13B,32'hB1490F62,32'hB08B6555,
    32'hBBD72268,32'hBA15485F,32'hB853F606,32'hB9919C31,32'hBCDE8AB4,32'hBD1CE083,32'hBF5A5EDA,32'hBE9834ED};

 logic [31:0] crctable3[256]= {32'h00000000,32'hB8BC6765,32'hAA09C88B,32'h12B5AFEE,32'h8F629757,32'h37DEF032,32'h256B5FDC,32'h9DD738B9,
    32'hC5B428EF,32'h7D084F8A,32'h6FBDE064,32'hD7018701,32'h4AD6BFB8,32'hF26AD8DD,32'hE0DF7733,32'h58631056,
    32'h5019579F,32'hE8A530FA,32'hFA109F14,32'h42ACF871,32'hDF7BC0C8,32'h67C7A7AD,32'h75720843,32'hCDCE6F26,
    32'h95AD7F70,32'h2D111815,32'h3FA4B7FB,32'h8718D09E,32'h1ACFE827,32'hA2738F42,32'hB0C620AC,32'h087A47C9,
    32'hA032AF3E,32'h188EC85B,32'h0A3B67B5,32'hB28700D0,32'h2F503869,32'h97EC5F0C,32'h8559F0E2,32'h3DE59787,
    32'h658687D1,32'hDD3AE0B4,32'hCF8F4F5A,32'h7733283F,32'hEAE41086,32'h525877E3,32'h40EDD80D,32'hF851BF68,
    32'hF02BF8A1,32'h48979FC4,32'h5A22302A,32'hE29E574F,32'h7F496FF6,32'hC7F50893,32'hD540A77D,32'h6DFCC018,
    32'h359FD04E,32'h8D23B72B,32'h9F9618C5,32'h272A7FA0,32'hBAFD4719,32'h0241207C,32'h10F48F92,32'hA848E8F7,
    32'h9B14583D,32'h23A83F58,32'h311D90B6,32'h89A1F7D3,32'h1476CF6A,32'hACCAA80F,32'hBE7F07E1,32'h06C36084,
    32'h5EA070D2,32'hE61C17B7,32'hF4A9B859,32'h4C15DF3C,32'hD1C2E785,32'h697E80E0,32'h7BCB2F0E,32'hC377486B,
    32'hCB0D0FA2,32'h73B168C7,32'h6104C729,32'hD9B8A04C,32'h446F98F5,32'hFCD3FF90,32'hEE66507E,32'h56DA371B,
    32'h0EB9274D,32'hB6054028,32'hA4B0EFC6,32'h1C0C88A3,32'h81DBB01A,32'h3967D77F,32'h2BD27891,32'h936E1FF4,
    32'h3B26F703,32'h839A9066,32'h912F3F88,32'h299358ED,32'hB4446054,32'h0CF80731,32'h1E4DA8DF,32'hA6F1CFBA,
    32'hFE92DFEC,32'h462EB889,32'h549B1767,32'hEC277002,32'h71F048BB,32'hC94C2FDE,32'hDBF98030,32'h6345E755,
    32'h6B3FA09C,32'hD383C7F9,32'hC1366817,32'h798A0F72,32'hE45D37CB,32'h5CE150AE,32'h4E54FF40,32'hF6E89825,
    32'hAE8B8873,32'h1637EF16,32'h048240F8,32'hBC3E279D,32'h21E91F24,32'h99557841,32'h8BE0D7AF,32'h335CB0CA,
    32'hED59B63B,32'h55E5D15E,32'h47507EB0,32'hFFEC19D5,32'h623B216C,32'hDA874609,32'hC832E9E7,32'h708E8E82,
    32'h28ED9ED4,32'h9051F9B1,32'h82E4565F,32'h3A58313A,32'hA78F0983,32'h1F336EE6,32'h0D86C108,32'hB53AA66D,
    32'hBD40E1A4,32'h05FC86C1,32'h1749292F,32'hAFF54E4A,32'h322276F3,32'h8A9E1196,32'h982BBE78,32'h2097D91D,
    32'h78F4C94B,32'hC048AE2E,32'hD2FD01C0,32'h6A4166A5,32'hF7965E1C,32'h4F2A3979,32'h5D9F9697,32'hE523F1F2,
    32'h4D6B1905,32'hF5D77E60,32'hE762D18E,32'h5FDEB6EB,32'hC2098E52,32'h7AB5E937,32'h680046D9,32'hD0BC21BC,
    32'h88DF31EA,32'h3063568F,32'h22D6F961,32'h9A6A9E04,32'h07BDA6BD,32'hBF01C1D8,32'hADB46E36,32'h15080953,
    32'h1D724E9A,32'hA5CE29FF,32'hB77B8611,32'h0FC7E174,32'h9210D9CD,32'h2AACBEA8,32'h38191146,32'h80A57623,
    32'hD8C66675,32'h607A0110,32'h72CFAEFE,32'hCA73C99B,32'h57A4F122,32'hEF189647,32'hFDAD39A9,32'h45115ECC,
    32'h764DEE06,32'hCEF18963,32'hDC44268D,32'h64F841E8,32'hF92F7951,32'h41931E34,32'h5326B1DA,32'hEB9AD6BF,
    32'hB3F9C6E9,32'h0B45A18C,32'h19F00E62,32'hA14C6907,32'h3C9B51BE,32'h842736DB,32'h96929935,32'h2E2EFE50,
    32'h2654B999,32'h9EE8DEFC,32'h8C5D7112,32'h34E11677,32'hA9362ECE,32'h118A49AB,32'h033FE645,32'hBB838120,
    32'hE3E09176,32'h5B5CF613,32'h49E959FD,32'hF1553E98,32'h6C820621,32'hD43E6144,32'hC68BCEAA,32'h7E37A9CF,
    32'hD67F4138,32'h6EC3265D,32'h7C7689B3,32'hC4CAEED6,32'h591DD66F,32'hE1A1B10A,32'hF3141EE4,32'h4BA87981,
    32'h13CB69D7,32'hAB770EB2,32'hB9C2A15C,32'h017EC639,32'h9CA9FE80,32'h241599E5,32'h36A0360B,32'h8E1C516E,
    32'h866616A7,32'h3EDA71C2,32'h2C6FDE2C,32'h94D3B949,32'h090481F0,32'hB1B8E695,32'hA30D497B,32'h1BB12E1E,
    32'h43D23E48,32'hFB6E592D,32'hE9DBF6C3,32'h516791A6,32'hCCB0A91F,32'h740CCE7A,32'h66B96194,32'hDE0506F1};
    
    logic [31:0] crctable4[256]={ 32'h00000000,32'h3D6029B0,32'h7AC05360,32'h47A07AD0,32'hF580A6C0,32'hC8E08F70,32'h8F40F5A0,32'hB220DC10,
    32'h30704BC1,32'h0D106271,32'h4AB018A1,32'h77D03111,32'hC5F0ED01,32'hF890C4B1,32'hBF30BE61,32'h825097D1,
    32'h60E09782,32'h5D80BE32,32'h1A20C4E2,32'h2740ED52,32'h95603142,32'hA80018F2,32'hEFA06222,32'hD2C04B92,
    32'h5090DC43,32'h6DF0F5F3,32'h2A508F23,32'h1730A693,32'hA5107A83,32'h98705333,32'hDFD029E3,32'hE2B00053,
    32'hC1C12F04,32'hFCA106B4,32'hBB017C64,32'h866155D4,32'h344189C4,32'h0921A074,32'h4E81DAA4,32'h73E1F314,
    32'hF1B164C5,32'hCCD14D75,32'h8B7137A5,32'hB6111E15,32'h0431C205,32'h3951EBB5,32'h7EF19165,32'h4391B8D5,
    32'hA121B886,32'h9C419136,32'hDBE1EBE6,32'hE681C256,32'h54A11E46,32'h69C137F6,32'h2E614D26,32'h13016496,
    32'h9151F347,32'hAC31DAF7,32'hEB91A027,32'hD6F18997,32'h64D15587,32'h59B17C37,32'h1E1106E7,32'h23712F57,
    32'h58F35849,32'h659371F9,32'h22330B29,32'h1F532299,32'hAD73FE89,32'h9013D739,32'hD7B3ADE9,32'hEAD38459,
    32'h68831388,32'h55E33A38,32'h124340E8,32'h2F236958,32'h9D03B548,32'hA0639CF8,32'hE7C3E628,32'hDAA3CF98,
    32'h3813CFCB,32'h0573E67B,32'h42D39CAB,32'h7FB3B51B,32'hCD93690B,32'hF0F340BB,32'hB7533A6B,32'h8A3313DB,
    32'h0863840A,32'h3503ADBA,32'h72A3D76A,32'h4FC3FEDA,32'hFDE322CA,32'hC0830B7A,32'h872371AA,32'hBA43581A,
    32'h9932774D,32'hA4525EFD,32'hE3F2242D,32'hDE920D9D,32'h6CB2D18D,32'h51D2F83D,32'h167282ED,32'h2B12AB5D,
    32'hA9423C8C,32'h9422153C,32'hD3826FEC,32'hEEE2465C,32'h5CC29A4C,32'h61A2B3FC,32'h2602C92C,32'h1B62E09C,
    32'hF9D2E0CF,32'hC4B2C97F,32'h8312B3AF,32'hBE729A1F,32'h0C52460F,32'h31326FBF,32'h7692156F,32'h4BF23CDF,
    32'hC9A2AB0E,32'hF4C282BE,32'hB362F86E,32'h8E02D1DE,32'h3C220DCE,32'h0142247E,32'h46E25EAE,32'h7B82771E,
    32'hB1E6B092,32'h8C869922,32'hCB26E3F2,32'hF646CA42,32'h44661652,32'h79063FE2,32'h3EA64532,32'h03C66C82,
    32'h8196FB53,32'hBCF6D2E3,32'hFB56A833,32'hC6368183,32'h74165D93,32'h49767423,32'h0ED60EF3,32'h33B62743,
    32'hD1062710,32'hEC660EA0,32'hABC67470,32'h96A65DC0,32'h248681D0,32'h19E6A860,32'h5E46D2B0,32'h6326FB00,
    32'hE1766CD1,32'hDC164561,32'h9BB63FB1,32'hA6D61601,32'h14F6CA11,32'h2996E3A1,32'h6E369971,32'h5356B0C1,
    32'h70279F96,32'h4D47B626,32'h0AE7CCF6,32'h3787E546,32'h85A73956,32'hB8C710E6,32'hFF676A36,32'hC2074386,
    32'h4057D457,32'h7D37FDE7,32'h3A978737,32'h07F7AE87,32'hB5D77297,32'h88B75B27,32'hCF1721F7,32'hF2770847,
    32'h10C70814,32'h2DA721A4,32'h6A075B74,32'h576772C4,32'hE547AED4,32'hD8278764,32'h9F87FDB4,32'hA2E7D404,
    32'h20B743D5,32'h1DD76A65,32'h5A7710B5,32'h67173905,32'hD537E515,32'hE857CCA5,32'hAFF7B675,32'h92979FC5,
    32'hE915E8DB,32'hD475C16B,32'h93D5BBBB,32'hAEB5920B,32'h1C954E1B,32'h21F567AB,32'h66551D7B,32'h5B3534CB,
    32'hD965A31A,32'hE4058AAA,32'hA3A5F07A,32'h9EC5D9CA,32'h2CE505DA,32'h11852C6A,32'h562556BA,32'h6B457F0A,
    32'h89F57F59,32'hB49556E9,32'hF3352C39,32'hCE550589,32'h7C75D999,32'h4115F029,32'h06B58AF9,32'h3BD5A349,
    32'hB9853498,32'h84E51D28,32'hC34567F8,32'hFE254E48,32'h4C059258,32'h7165BBE8,32'h36C5C138,32'h0BA5E888,
    32'h28D4C7DF,32'h15B4EE6F,32'h521494BF,32'h6F74BD0F,32'hDD54611F,32'hE03448AF,32'hA794327F,32'h9AF41BCF,
    32'h18A48C1E,32'h25C4A5AE,32'h6264DF7E,32'h5F04F6CE,32'hED242ADE,32'hD044036E,32'h97E479BE,32'hAA84500E,
    32'h4834505D,32'h755479ED,32'h32F4033D,32'h0F942A8D,32'hBDB4F69D,32'h80D4DF2D,32'hC774A5FD,32'hFA148C4D,
    32'h78441B9C,32'h4524322C,32'h028448FC,32'h3FE4614C,32'h8DC4BD5C,32'hB0A494EC,32'hF704EE3C,32'hCA64C78C};
    
    logic [31:0] crctable5[256]={32'h00000000,32'hCB5CD3A5,32'h4DC8A10B,32'h869472AE,32'h9B914216,32'h50CD91B3,32'hD659E31D,32'h1D0530B8,
    32'hEC53826D,32'h270F51C8,32'hA19B2366,32'h6AC7F0C3,32'h77C2C07B,32'hBC9E13DE,32'h3A0A6170,32'hF156B2D5,
    32'h03D6029B,32'hC88AD13E,32'h4E1EA390,32'h85427035,32'h9847408D,32'h531B9328,32'hD58FE186,32'h1ED33223,
    32'hEF8580F6,32'h24D95353,32'hA24D21FD,32'h6911F258,32'h7414C2E0,32'hBF481145,32'h39DC63EB,32'hF280B04E,
    32'h07AC0536,32'hCCF0D693,32'h4A64A43D,32'h81387798,32'h9C3D4720,32'h57619485,32'hD1F5E62B,32'h1AA9358E,
    32'hEBFF875B,32'h20A354FE,32'hA6372650,32'h6D6BF5F5,32'h706EC54D,32'hBB3216E8,32'h3DA66446,32'hF6FAB7E3,
    32'h047A07AD,32'hCF26D408,32'h49B2A6A6,32'h82EE7503,32'h9FEB45BB,32'h54B7961E,32'hD223E4B0,32'h197F3715,
    32'hE82985C0,32'h23755665,32'hA5E124CB,32'h6EBDF76E,32'h73B8C7D6,32'hB8E41473,32'h3E7066DD,32'hF52CB578,
    32'h0F580A6C,32'hC404D9C9,32'h4290AB67,32'h89CC78C2,32'h94C9487A,32'h5F959BDF,32'hD901E971,32'h125D3AD4,
    32'hE30B8801,32'h28575BA4,32'hAEC3290A,32'h659FFAAF,32'h789ACA17,32'hB3C619B2,32'h35526B1C,32'hFE0EB8B9,
    32'h0C8E08F7,32'hC7D2DB52,32'h4146A9FC,32'h8A1A7A59,32'h971F4AE1,32'h5C439944,32'hDAD7EBEA,32'h118B384F,
    32'hE0DD8A9A,32'h2B81593F,32'hAD152B91,32'h6649F834,32'h7B4CC88C,32'hB0101B29,32'h36846987,32'hFDD8BA22,
    32'h08F40F5A,32'hC3A8DCFF,32'h453CAE51,32'h8E607DF4,32'h93654D4C,32'h58399EE9,32'hDEADEC47,32'h15F13FE2,
    32'hE4A78D37,32'h2FFB5E92,32'hA96F2C3C,32'h6233FF99,32'h7F36CF21,32'hB46A1C84,32'h32FE6E2A,32'hF9A2BD8F,
    32'h0B220DC1,32'hC07EDE64,32'h46EAACCA,32'h8DB67F6F,32'h90B34FD7,32'h5BEF9C72,32'hDD7BEEDC,32'h16273D79,
    32'hE7718FAC,32'h2C2D5C09,32'hAAB92EA7,32'h61E5FD02,32'h7CE0CDBA,32'hB7BC1E1F,32'h31286CB1,32'hFA74BF14,
    32'h1EB014D8,32'hD5ECC77D,32'h5378B5D3,32'h98246676,32'h852156CE,32'h4E7D856B,32'hC8E9F7C5,32'h03B52460,
    32'hF2E396B5,32'h39BF4510,32'hBF2B37BE,32'h7477E41B,32'h6972D4A3,32'hA22E0706,32'h24BA75A8,32'hEFE6A60D,
    32'h1D661643,32'hD63AC5E6,32'h50AEB748,32'h9BF264ED,32'h86F75455,32'h4DAB87F0,32'hCB3FF55E,32'h006326FB,
    32'hF135942E,32'h3A69478B,32'hBCFD3525,32'h77A1E680,32'h6AA4D638,32'hA1F8059D,32'h276C7733,32'hEC30A496,
    32'h191C11EE,32'hD240C24B,32'h54D4B0E5,32'h9F886340,32'h828D53F8,32'h49D1805D,32'hCF45F2F3,32'h04192156,
    32'hF54F9383,32'h3E134026,32'hB8873288,32'h73DBE12D,32'h6EDED195,32'hA5820230,32'h2316709E,32'hE84AA33B,
    32'h1ACA1375,32'hD196C0D0,32'h5702B27E,32'h9C5E61DB,32'h815B5163,32'h4A0782C6,32'hCC93F068,32'h07CF23CD,
    32'hF6999118,32'h3DC542BD,32'hBB513013,32'h700DE3B6,32'h6D08D30E,32'hA65400AB,32'h20C07205,32'hEB9CA1A0,
    32'h11E81EB4,32'hDAB4CD11,32'h5C20BFBF,32'h977C6C1A,32'h8A795CA2,32'h41258F07,32'hC7B1FDA9,32'h0CED2E0C,
    32'hFDBB9CD9,32'h36E74F7C,32'hB0733DD2,32'h7B2FEE77,32'h662ADECF,32'hAD760D6A,32'h2BE27FC4,32'hE0BEAC61,
    32'h123E1C2F,32'hD962CF8A,32'h5FF6BD24,32'h94AA6E81,32'h89AF5E39,32'h42F38D9C,32'hC467FF32,32'h0F3B2C97,
    32'hFE6D9E42,32'h35314DE7,32'hB3A53F49,32'h78F9ECEC,32'h65FCDC54,32'hAEA00FF1,32'h28347D5F,32'hE368AEFA,
    32'h16441B82,32'hDD18C827,32'h5B8CBA89,32'h90D0692C,32'h8DD55994,32'h46898A31,32'hC01DF89F,32'h0B412B3A,
    32'hFA1799EF,32'h314B4A4A,32'hB7DF38E4,32'h7C83EB41,32'h6186DBF9,32'hAADA085C,32'h2C4E7AF2,32'hE712A957,
    32'h15921919,32'hDECECABC,32'h585AB812,32'h93066BB7,32'h8E035B0F,32'h455F88AA,32'hC3CBFA04,32'h089729A1,
    32'hF9C19B74,32'h329D48D1,32'hB4093A7F,32'h7F55E9DA,32'h6250D962,32'hA90C0AC7,32'h2F987869,32'hE4C4ABCC};
    
  logic [31:0] crctable6[256]= {32'h00000000,32'hA6770BB4,32'h979F1129,32'h31E81A9D,32'hF44F2413,32'h52382FA7,32'h63D0353A,32'hC5A73E8E,
    32'h33EF4E67,32'h959845D3,32'hA4705F4E,32'h020754FA,32'hC7A06A74,32'h61D761C0,32'h503F7B5D,32'hF64870E9,
    32'h67DE9CCE,32'hC1A9977A,32'hF0418DE7,32'h56368653,32'h9391B8DD,32'h35E6B369,32'h040EA9F4,32'hA279A240,
    32'h5431D2A9,32'hF246D91D,32'hC3AEC380,32'h65D9C834,32'hA07EF6BA,32'h0609FD0E,32'h37E1E793,32'h9196EC27,
    32'hCFBD399C,32'h69CA3228,32'h582228B5,32'hFE552301,32'h3BF21D8F,32'h9D85163B,32'hAC6D0CA6,32'h0A1A0712,
    32'hFC5277FB,32'h5A257C4F,32'h6BCD66D2,32'hCDBA6D66,32'h081D53E8,32'hAE6A585C,32'h9F8242C1,32'h39F54975,
    32'hA863A552,32'h0E14AEE6,32'h3FFCB47B,32'h998BBFCF,32'h5C2C8141,32'hFA5B8AF5,32'hCBB39068,32'h6DC49BDC,
    32'h9B8CEB35,32'h3DFBE081,32'h0C13FA1C,32'hAA64F1A8,32'h6FC3CF26,32'hC9B4C492,32'hF85CDE0F,32'h5E2BD5BB,
    32'h440B7579,32'hE27C7ECD,32'hD3946450,32'h75E36FE4,32'hB044516A,32'h16335ADE,32'h27DB4043,32'h81AC4BF7,
    32'h77E43B1E,32'hD19330AA,32'hE07B2A37,32'h460C2183,32'h83AB1F0D,32'h25DC14B9,32'h14340E24,32'hB2430590,
    32'h23D5E9B7,32'h85A2E203,32'hB44AF89E,32'h123DF32A,32'hD79ACDA4,32'h71EDC610,32'h4005DC8D,32'hE672D739,
    32'h103AA7D0,32'hB64DAC64,32'h87A5B6F9,32'h21D2BD4D,32'hE47583C3,32'h42028877,32'h73EA92EA,32'hD59D995E,
    32'h8BB64CE5,32'h2DC14751,32'h1C295DCC,32'hBA5E5678,32'h7FF968F6,32'hD98E6342,32'hE86679DF,32'h4E11726B,
    32'hB8590282,32'h1E2E0936,32'h2FC613AB,32'h89B1181F,32'h4C162691,32'hEA612D25,32'hDB8937B8,32'h7DFE3C0C,
    32'hEC68D02B,32'h4A1FDB9F,32'h7BF7C102,32'hDD80CAB6,32'h1827F438,32'hBE50FF8C,32'h8FB8E511,32'h29CFEEA5,
    32'hDF879E4C,32'h79F095F8,32'h48188F65,32'hEE6F84D1,32'h2BC8BA5F,32'h8DBFB1EB,32'hBC57AB76,32'h1A20A0C2,
    32'h8816EAF2,32'h2E61E146,32'h1F89FBDB,32'hB9FEF06F,32'h7C59CEE1,32'hDA2EC555,32'hEBC6DFC8,32'h4DB1D47C,
    32'hBBF9A495,32'h1D8EAF21,32'h2C66B5BC,32'h8A11BE08,32'h4FB68086,32'hE9C18B32,32'hD82991AF,32'h7E5E9A1B,
    32'hEFC8763C,32'h49BF7D88,32'h78576715,32'hDE206CA1,32'h1B87522F,32'hBDF0599B,32'h8C184306,32'h2A6F48B2,
    32'hDC27385B,32'h7A5033EF,32'h4BB82972,32'hEDCF22C6,32'h28681C48,32'h8E1F17FC,32'hBFF70D61,32'h198006D5,
    32'h47ABD36E,32'hE1DCD8DA,32'hD034C247,32'h7643C9F3,32'hB3E4F77D,32'h1593FCC9,32'h247BE654,32'h820CEDE0,
    32'h74449D09,32'hD23396BD,32'hE3DB8C20,32'h45AC8794,32'h800BB91A,32'h267CB2AE,32'h1794A833,32'hB1E3A387,
    32'h20754FA0,32'h86024414,32'hB7EA5E89,32'h119D553D,32'hD43A6BB3,32'h724D6007,32'h43A57A9A,32'hE5D2712E,
    32'h139A01C7,32'hB5ED0A73,32'h840510EE,32'h22721B5A,32'hE7D525D4,32'h41A22E60,32'h704A34FD,32'hD63D3F49,
    32'hCC1D9F8B,32'h6A6A943F,32'h5B828EA2,32'hFDF58516,32'h3852BB98,32'h9E25B02C,32'hAFCDAAB1,32'h09BAA105,
    32'hFFF2D1EC,32'h5985DA58,32'h686DC0C5,32'hCE1ACB71,32'h0BBDF5FF,32'hADCAFE4B,32'h9C22E4D6,32'h3A55EF62,
    32'hABC30345,32'h0DB408F1,32'h3C5C126C,32'h9A2B19D8,32'h5F8C2756,32'hF9FB2CE2,32'hC813367F,32'h6E643DCB,
    32'h982C4D22,32'h3E5B4696,32'h0FB35C0B,32'hA9C457BF,32'h6C636931,32'hCA146285,32'hFBFC7818,32'h5D8B73AC,
    32'h03A0A617,32'hA5D7ADA3,32'h943FB73E,32'h3248BC8A,32'hF7EF8204,32'h519889B0,32'h6070932D,32'hC6079899,
    32'h304FE870,32'h9638E3C4,32'hA7D0F959,32'h01A7F2ED,32'hC400CC63,32'h6277C7D7,32'h539FDD4A,32'hF5E8D6FE,
    32'h647E3AD9,32'hC209316D,32'hF3E12BF0,32'h55962044,32'h90311ECA,32'h3646157E,32'h07AE0FE3,32'hA1D90457,
    32'h579174BE,32'hF1E67F0A,32'hC00E6597,32'h66796E23,32'hA3DE50AD,32'h05A95B19,32'h34414184,32'h92364A30};
    
    logic [31:0] crctable7[256]={32'h00000000,32'hCCAA009E,32'h4225077D,32'h8E8F07E3,32'h844A0EFA,32'h48E00E64,32'hC66F0987,32'h0AC50919,
    32'hD3E51BB5,32'h1F4F1B2B,32'h91C01CC8,32'h5D6A1C56,32'h57AF154F,32'h9B0515D1,32'h158A1232,32'hD92012AC,
    32'h7CBB312B,32'hB01131B5,32'h3E9E3656,32'hF23436C8,32'hF8F13FD1,32'h345B3F4F,32'hBAD438AC,32'h767E3832,
    32'hAF5E2A9E,32'h63F42A00,32'hED7B2DE3,32'h21D12D7D,32'h2B142464,32'hE7BE24FA,32'h69312319,32'hA59B2387,
    32'hF9766256,32'h35DC62C8,32'hBB53652B,32'h77F965B5,32'h7D3C6CAC,32'hB1966C32,32'h3F196BD1,32'hF3B36B4F,
    32'h2A9379E3,32'hE639797D,32'h68B67E9E,32'hA41C7E00,32'hAED97719,32'h62737787,32'hECFC7064,32'h205670FA,
    32'h85CD537D,32'h496753E3,32'hC7E85400,32'h0B42549E,32'h01875D87,32'hCD2D5D19,32'h43A25AFA,32'h8F085A64,
    32'h562848C8,32'h9A824856,32'h140D4FB5,32'hD8A74F2B,32'hD2624632,32'h1EC846AC,32'h9047414F,32'h5CED41D1,
    32'h299DC2ED,32'hE537C273,32'h6BB8C590,32'hA712C50E,32'hADD7CC17,32'h617DCC89,32'hEFF2CB6A,32'h2358CBF4,
    32'hFA78D958,32'h36D2D9C6,32'hB85DDE25,32'h74F7DEBB,32'h7E32D7A2,32'hB298D73C,32'h3C17D0DF,32'hF0BDD041,
    32'h5526F3C6,32'h998CF358,32'h1703F4BB,32'hDBA9F425,32'hD16CFD3C,32'h1DC6FDA2,32'h9349FA41,32'h5FE3FADF,
    32'h86C3E873,32'h4A69E8ED,32'hC4E6EF0E,32'h084CEF90,32'h0289E689,32'hCE23E617,32'h40ACE1F4,32'h8C06E16A,
    32'hD0EBA0BB,32'h1C41A025,32'h92CEA7C6,32'h5E64A758,32'h54A1AE41,32'h980BAEDF,32'h1684A93C,32'hDA2EA9A2,
    32'h030EBB0E,32'hCFA4BB90,32'h412BBC73,32'h8D81BCED,32'h8744B5F4,32'h4BEEB56A,32'hC561B289,32'h09CBB217,
    32'hAC509190,32'h60FA910E,32'hEE7596ED,32'h22DF9673,32'h281A9F6A,32'hE4B09FF4,32'h6A3F9817,32'hA6959889,
    32'h7FB58A25,32'hB31F8ABB,32'h3D908D58,32'hF13A8DC6,32'hFBFF84DF,32'h37558441,32'hB9DA83A2,32'h7570833C,
    32'h533B85DA,32'h9F918544,32'h111E82A7,32'hDDB48239,32'hD7718B20,32'h1BDB8BBE,32'h95548C5D,32'h59FE8CC3,
    32'h80DE9E6F,32'h4C749EF1,32'hC2FB9912,32'h0E51998C,32'h04949095,32'hC83E900B,32'h46B197E8,32'h8A1B9776,
    32'h2F80B4F1,32'hE32AB46F,32'h6DA5B38C,32'hA10FB312,32'hABCABA0B,32'h6760BA95,32'hE9EFBD76,32'h2545BDE8,
    32'hFC65AF44,32'h30CFAFDA,32'hBE40A839,32'h72EAA8A7,32'h782FA1BE,32'hB485A120,32'h3A0AA6C3,32'hF6A0A65D,
    32'hAA4DE78C,32'h66E7E712,32'hE868E0F1,32'h24C2E06F,32'h2E07E976,32'hE2ADE9E8,32'h6C22EE0B,32'hA088EE95,
    32'h79A8FC39,32'hB502FCA7,32'h3B8DFB44,32'hF727FBDA,32'hFDE2F2C3,32'h3148F25D,32'hBFC7F5BE,32'h736DF520,
    32'hD6F6D6A7,32'h1A5CD639,32'h94D3D1DA,32'h5879D144,32'h52BCD85D,32'h9E16D8C3,32'h1099DF20,32'hDC33DFBE,
    32'h0513CD12,32'hC9B9CD8C,32'h4736CA6F,32'h8B9CCAF1,32'h8159C3E8,32'h4DF3C376,32'hC37CC495,32'h0FD6C40B,
    32'h7AA64737,32'hB60C47A9,32'h3883404A,32'hF42940D4,32'hFEEC49CD,32'h32464953,32'hBCC94EB0,32'h70634E2E,
    32'hA9435C82,32'h65E95C1C,32'hEB665BFF,32'h27CC5B61,32'h2D095278,32'hE1A352E6,32'h6F2C5505,32'hA386559B,
    32'h061D761C,32'hCAB77682,32'h44387161,32'h889271FF,32'h825778E6,32'h4EFD7878,32'hC0727F9B,32'h0CD87F05,
    32'hD5F86DA9,32'h19526D37,32'h97DD6AD4,32'h5B776A4A,32'h51B26353,32'h9D1863CD,32'h1397642E,32'hDF3D64B0,
    32'h83D02561,32'h4F7A25FF,32'hC1F5221C,32'h0D5F2282,32'h079A2B9B,32'hCB302B05,32'h45BF2CE6,32'h89152C78,
    32'h50353ED4,32'h9C9F3E4A,32'h121039A9,32'hDEBA3937,32'hD47F302E,32'h18D530B0,32'h965A3753,32'h5AF037CD,
    32'hFF6B144A,32'h33C114D4,32'hBD4E1337,32'h71E413A9,32'h7B211AB0,32'hB78B1A2E,32'h39041DCD,32'hF5AE1D53,
    32'h2C8E0FFF,32'hE0240F61,32'h6EAB0882,32'hA201081C,32'hA8C40105,32'h646E019B,32'hEAE10678,32'h264B06E6};
    
    
    
    
    logic  [31:0]crc_d[10:0];
    logic  [31:0]crc_q;
    logic  [31:0]my_crc;
    
    always_comb begin
    crc_d[0]  = ~old_crc_i;
    crc_d[1]  = crc_d[0]^ data_i[63:32]; 
    crc_d[2]  = crctable4[crc_d[1][7:0]];
    crc_d[3]  = crctable5[crc_d[1][15:8]];
    crc_d[4]  = crctable6[crc_d[1][23:16]];
    crc_d[5]  = crctable7[crc_d[1][31:24]];
   // my_crc = 32'h47eaa88b;
    crc_d[6]  = crctable0[data_i[7:0]  ];
    crc_d[7]  = crctable1[data_i[15:8] ];
    crc_d[8]  = crctable2[data_i[23:16]];
    crc_d[9]  = crctable3[data_i[31:24]];
    crc_d[10] = crc_d[2]^crc_d[3]^ crc_d[4]^crc_d[5]^crc_d[6]^crc_d[7]^ crc_d[8]^crc_d[9];      
    end       
     /*always_ff @(posedge clk_i or negedge rst_i) begin 
        if (rst_i ==1'b0) begin
                crc_q       <=  0;
        end
        else 
                crc_q        <= crc_d;
        end*/
    assign new_crc_o = ~crc_d[10];
endmodule
